module reg_16 (
    
);
    
endmodule